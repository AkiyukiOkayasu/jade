.title KiCad schematic
J8 GND GND Net-_J8-Pad3_ PJ302M
C1 +12V GND 10u
J1 GND GND Net-_J1-Pad3_ PJ302M
Q1 Net-_D1-Pad1_ GND /GATE_IN1 MMBT3904
R1 Net-_D1-Pad1_ Net-_J1-Pad3_ 100k
R5 GND Net-_D1-Pad1_ 100k
J2 GND GND Net-_J2-Pad3_ PJ302M
Q2 Net-_D2-Pad1_ GND /GATE_IN2 MMBT3904
R2 Net-_D2-Pad1_ Net-_J2-Pad3_ 100k
R6 GND Net-_D2-Pad1_ 100k
J3 GND GND Net-_J3-Pad3_ PJ302M
Q3 Net-_D3-Pad1_ GND /GATE_IN3 MMBT3904
R3 Net-_D3-Pad1_ Net-_J3-Pad3_ 100k
R7 GND Net-_D3-Pad1_ 100k
J4 GND GND Net-_J4-Pad3_ PJ302M
Q4 Net-_D4-Pad1_ GND /GATE_IN4 MMBT3904
R4 Net-_D4-Pad1_ Net-_J4-Pad3_ 100k
R8 GND Net-_D4-Pad1_ 100k
U2 Net-_R14-Pad1_ Net-_R11-Pad1_ Net-_R12-Pad1_ GND Net-_R10-Pad1_ Net-_R13-Pad2_ Net-_R13-Pad1_ +12V LM358
R12 Net-_R12-Pad1_ /CLOCK_OUT 10k
R11 Net-_R11-Pad1_ GND 39k
R14 Net-_R14-Pad1_ Net-_R11-Pad1_ 56k
R16 Net-_J8-Pad3_ Net-_R14-Pad1_ 1k
J7 GND GND Net-_J7-Pad3_ PJ302M
R10 Net-_R10-Pad1_ /GATE_OUT 10k
R9 Net-_R13-Pad2_ GND 39k
R13 Net-_R13-Pad1_ Net-_R13-Pad2_ 56k
R15 Net-_J7-Pad3_ Net-_R13-Pad1_ 1k
J5 Net-_D5-Pad2_ Net-_D5-Pad2_ GND GND GND GND GND GND NC_01 NC_02 Conn_02x05_Odd_Even
D5 +12V Net-_D5-Pad2_ 1N5819HW
C2 +12V GND 0.1u
U1 NC_03 NC_04 /CLOCK_OUT /GATE_OUT /SDA /SCL /GATE_IN1 NC_05 /GATE_IN2 /GATE_IN3 /GATE_IN4 NC_06 GND NC_07 NC_08 GND NC_09 NC_10 NC_11 GND SeeeduinoXIAO
J6 /SDA /SDA /SCL /SCL GND GND Conn_02x03_Odd_Even
D4 Net-_D4-Pad1_ GND 1N4148W
D1 Net-_D1-Pad1_ GND 1N4148W
D2 Net-_D2-Pad1_ GND 1N4148W
D3 Net-_D3-Pad1_ GND 1N4148W
.end
